-- Name:				division.vhd
-- Filetype:		VHDL Testbench
-- Date:				23 september 2019
-- Description:	psuedo-divides tix to calculate RPM
-- Author:			Bjoern van Rozelaar for PRODIG-PETERS-PG1
-- State:			Testing
-- Error:			-
-- Version:			1.0

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--Empty entity
entity tb_division is
end entity

--The architecture
architecture sim of tb_division is
	port
	(
	
	)
	;
end component tb_division;

--Signalen om te monitoren


--S