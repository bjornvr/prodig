-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Sep 18 13:33:55 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY RPM_CLOCK IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Hallsensor : IN STD_LOGIC := '0';
        Start_count : OUT STD_LOGIC
    );
END RPM_CLOCK;

ARCHITECTURE BEHAVIOR OF RPM_CLOCK IS
    TYPE type_fstate IS (invalide,start_count,calculate,compair,start);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='0') THEN
            fstate <= start;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,Hallsensor)
    BEGIN
        Start_count <= '0';
        CASE fstate IS
            WHEN invalide =>
                reg_fstate <= start;
            WHEN start_count =>
                IF (NOT((Hallsensor = '1'))) THEN
                    reg_fstate <= compair;
                ELSIF ((Hallsensor = '1')) THEN
                    reg_fstate <= start_count;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= start_count;
                END IF;

                Start_count <= '1';
            WHEN calculate =>
                reg_fstate <= start;

                Start_count <= '0';
            WHEN compair =>
                IF ((Hallsensor = '1')) THEN
                    reg_fstate <= calculate;
                ELSIF (NOT((Hallsensor = '1'))) THEN
                    reg_fstate <= invalide;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= compair;
                END IF;
            WHEN start =>
                IF ((Hallsensor = '1')) THEN
                    reg_fstate <= start_count;
                ELSIF (NOT((Hallsensor = '1'))) THEN
                    reg_fstate <= start;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= start;
                END IF;

                Start_count <= '0';
            WHEN OTHERS => 
                Start_count <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
